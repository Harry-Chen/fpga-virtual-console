
module Probe (
	source,
	probe);	

	output	[15:0]	source;
	input	[127:0]	probe;
endmodule

module FpgaVirtualConsole(
input hello,
output world
);

assign world = hello;

endmodule
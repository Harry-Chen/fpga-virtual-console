module Color256Decoder(
	input  [7:0] code,
	output [8:0] color
);

always_comb
begin
	case(code)
		8'h00: color = 9'b000_000_000; // Black
		8'h01: color = 9'b100_000_000; // Maroon
		8'h02: color = 9'b000_100_000; // Green
		8'h03: color = 9'b100_100_000; // Olive
		8'h04: color = 9'b000_000_100; // Navy
		8'h05: color = 9'b100_000_100; // Purple
		8'h06: color = 9'b000_100_100; // Teal
		8'h07: color = 9'b110_110_110; // Silver
		8'h08: color = 9'b100_100_100; // Grey
		8'h09: color = 9'b111_000_000; // Red
		8'h0a: color = 9'b000_111_000; // Lime
		8'h0b: color = 9'b111_111_000; // Yellow
		8'h0c: color = 9'b000_000_111; // Blue
		8'h0d: color = 9'b111_000_111; // Fuchsia
		8'h0e: color = 9'b000_111_111; // Aqua
		8'h0f: color = 9'b111_111_111; // White
		8'h10: color = 9'b000_000_000; // Grey0
		8'h11: color = 9'b000_000_010; // NavyBlue
		8'h12: color = 9'b000_000_100; // DarkBlue
		8'h13: color = 9'b000_000_101; // Blue3
		8'h14: color = 9'b000_000_110; // Blue3
		8'h15: color = 9'b000_000_111; // Blue1
		8'h16: color = 9'b000_010_000; // DarkGreen
		8'h17: color = 9'b000_010_010; // DeepSkyBlue4
		8'h18: color = 9'b000_010_100; // DeepSkyBlue4
		8'h19: color = 9'b000_010_101; // DeepSkyBlue4
		8'h1a: color = 9'b000_010_110; // DodgerBlue3
		8'h1b: color = 9'b000_010_111; // DodgerBlue2
		8'h1c: color = 9'b000_100_000; // Green4
		8'h1d: color = 9'b000_100_010; // SpringGreen4
		8'h1e: color = 9'b000_100_100; // Turquoise4
		8'h1f: color = 9'b000_100_101; // DeepSkyBlue3
		8'h20: color = 9'b000_100_110; // DeepSkyBlue3
		8'h21: color = 9'b000_100_111; // DodgerBlue1
		8'h22: color = 9'b000_101_000; // Green3
		8'h23: color = 9'b000_101_010; // SpringGreen3
		8'h24: color = 9'b000_101_100; // DarkCyan
		8'h25: color = 9'b000_101_101; // LightSeaGreen
		8'h26: color = 9'b000_101_110; // DeepSkyBlue2
		8'h27: color = 9'b000_101_111; // DeepSkyBlue1
		8'h28: color = 9'b000_110_000; // Green3
		8'h29: color = 9'b000_110_010; // SpringGreen3
		8'h2a: color = 9'b000_110_100; // SpringGreen2
		8'h2b: color = 9'b000_110_101; // Cyan3
		8'h2c: color = 9'b000_110_110; // DarkTurquoise
		8'h2d: color = 9'b000_110_111; // Turquoise2
		8'h2e: color = 9'b000_111_000; // Green1
		8'h2f: color = 9'b000_111_010; // SpringGreen2
		8'h30: color = 9'b000_111_100; // SpringGreen1
		8'h31: color = 9'b000_111_101; // MediumSpringGreen
		8'h32: color = 9'b000_111_110; // Cyan2
		8'h33: color = 9'b000_111_111; // Cyan1
		8'h34: color = 9'b010_000_000; // DarkRed
		8'h35: color = 9'b010_000_010; // DeepPink4
		8'h36: color = 9'b010_000_100; // Purple4
		8'h37: color = 9'b010_000_101; // Purple4
		8'h38: color = 9'b010_000_110; // Purple3
		8'h39: color = 9'b010_000_111; // BlueViolet
		8'h3a: color = 9'b010_010_000; // Orange4
		8'h3b: color = 9'b010_010_010; // Grey37
		8'h3c: color = 9'b010_010_100; // MediumPurple4
		8'h3d: color = 9'b010_010_101; // SlateBlue3
		8'h3e: color = 9'b010_010_110; // SlateBlue3
		8'h3f: color = 9'b010_010_111; // RoyalBlue1
		8'h40: color = 9'b010_100_000; // Chartreuse4
		8'h41: color = 9'b010_100_010; // DarkSeaGreen4
		8'h42: color = 9'b010_100_100; // PaleTurquoise4
		8'h43: color = 9'b010_100_101; // SteelBlue
		8'h44: color = 9'b010_100_110; // SteelBlue3
		8'h45: color = 9'b010_100_111; // CornflowerBlue
		8'h46: color = 9'b010_101_000; // Chartreuse3
		8'h47: color = 9'b010_101_010; // DarkSeaGreen4
		8'h48: color = 9'b010_101_100; // CadetBlue
		8'h49: color = 9'b010_101_101; // CadetBlue
		8'h4a: color = 9'b010_101_110; // SkyBlue3
		8'h4b: color = 9'b010_101_111; // SteelBlue1
		8'h4c: color = 9'b010_110_000; // Chartreuse3
		8'h4d: color = 9'b010_110_010; // PaleGreen3
		8'h4e: color = 9'b010_110_100; // SeaGreen3
		8'h4f: color = 9'b010_110_101; // Aquamarine3
		8'h50: color = 9'b010_110_110; // MediumTurquoise
		8'h51: color = 9'b010_110_111; // SteelBlue1
		8'h52: color = 9'b010_111_000; // Chartreuse2
		8'h53: color = 9'b010_111_010; // SeaGreen2
		8'h54: color = 9'b010_111_100; // SeaGreen1
		8'h55: color = 9'b010_111_101; // SeaGreen1
		8'h56: color = 9'b010_111_110; // Aquamarine1
		8'h57: color = 9'b010_111_111; // DarkSlateGray2
		8'h58: color = 9'b100_000_000; // DarkRed
		8'h59: color = 9'b100_000_010; // DeepPink4
		8'h5a: color = 9'b100_000_100; // DarkMagenta
		8'h5b: color = 9'b100_000_101; // DarkMagenta
		8'h5c: color = 9'b100_000_110; // DarkViolet
		8'h5d: color = 9'b100_000_111; // Purple
		8'h5e: color = 9'b100_010_000; // Orange4
		8'h5f: color = 9'b100_010_010; // LightPink4
		8'h60: color = 9'b100_010_100; // Plum4
		8'h61: color = 9'b100_010_101; // MediumPurple3
		8'h62: color = 9'b100_010_110; // MediumPurple3
		8'h63: color = 9'b100_010_111; // SlateBlue1
		8'h64: color = 9'b100_100_000; // Yellow4
		8'h65: color = 9'b100_100_010; // Wheat4
		8'h66: color = 9'b100_100_100; // Grey53
		8'h67: color = 9'b100_100_101; // LightSlateGrey
		8'h68: color = 9'b100_100_110; // MediumPurple
		8'h69: color = 9'b100_100_111; // LightSlateBlue
		8'h6a: color = 9'b100_101_000; // Yellow4
		8'h6b: color = 9'b100_101_010; // DarkOliveGreen3
		8'h6c: color = 9'b100_101_100; // DarkSeaGreen
		8'h6d: color = 9'b100_101_101; // LightSkyBlue3
		8'h6e: color = 9'b100_101_110; // LightSkyBlue3
		8'h6f: color = 9'b100_101_111; // SkyBlue2
		8'h70: color = 9'b100_110_000; // Chartreuse2
		8'h71: color = 9'b100_110_010; // DarkOliveGreen3
		8'h72: color = 9'b100_110_100; // PaleGreen3
		8'h73: color = 9'b100_110_101; // DarkSeaGreen3
		8'h74: color = 9'b100_110_110; // DarkSlateGray3
		8'h75: color = 9'b100_110_111; // SkyBlue1
		8'h76: color = 9'b100_111_000; // Chartreuse1
		8'h77: color = 9'b100_111_010; // LightGreen
		8'h78: color = 9'b100_111_100; // LightGreen
		8'h79: color = 9'b100_111_101; // PaleGreen1
		8'h7a: color = 9'b100_111_110; // Aquamarine1
		8'h7b: color = 9'b100_111_111; // DarkSlateGray1
		8'h7c: color = 9'b101_000_000; // Red3
		8'h7d: color = 9'b101_000_010; // DeepPink4
		8'h7e: color = 9'b101_000_100; // MediumVioletRed
		8'h7f: color = 9'b101_000_101; // Magenta3
		8'h80: color = 9'b101_000_110; // DarkViolet
		8'h81: color = 9'b101_000_111; // Purple
		8'h82: color = 9'b101_010_000; // DarkOrange3
		8'h83: color = 9'b101_010_010; // IndianRed
		8'h84: color = 9'b101_010_100; // HotPink3
		8'h85: color = 9'b101_010_101; // MediumOrchid3
		8'h86: color = 9'b101_010_110; // MediumOrchid
		8'h87: color = 9'b101_010_111; // MediumPurple2
		8'h88: color = 9'b101_100_000; // DarkGoldenrod
		8'h89: color = 9'b101_100_010; // LightSalmon3
		8'h8a: color = 9'b101_100_100; // RosyBrown
		8'h8b: color = 9'b101_100_101; // Grey63
		8'h8c: color = 9'b101_100_110; // MediumPurple2
		8'h8d: color = 9'b101_100_111; // MediumPurple1
		8'h8e: color = 9'b101_101_000; // Gold3
		8'h8f: color = 9'b101_101_010; // DarkKhaki
		8'h90: color = 9'b101_101_100; // NavajoWhite3
		8'h91: color = 9'b101_101_101; // Grey69
		8'h92: color = 9'b101_101_110; // LightSteelBlue3
		8'h93: color = 9'b101_101_111; // LightSteelBlue
		8'h94: color = 9'b101_110_000; // Yellow3
		8'h95: color = 9'b101_110_010; // DarkOliveGreen3
		8'h96: color = 9'b101_110_100; // DarkSeaGreen3
		8'h97: color = 9'b101_110_101; // DarkSeaGreen2
		8'h98: color = 9'b101_110_110; // LightCyan3
		8'h99: color = 9'b101_110_111; // LightSkyBlue1
		8'h9a: color = 9'b101_111_000; // GreenYellow
		8'h9b: color = 9'b101_111_010; // DarkOliveGreen2
		8'h9c: color = 9'b101_111_100; // PaleGreen1
		8'h9d: color = 9'b101_111_101; // DarkSeaGreen2
		8'h9e: color = 9'b101_111_110; // DarkSeaGreen1
		8'h9f: color = 9'b101_111_111; // PaleTurquoise1
		8'ha0: color = 9'b110_000_000; // Red3
		8'ha1: color = 9'b110_000_010; // DeepPink3
		8'ha2: color = 9'b110_000_100; // DeepPink3
		8'ha3: color = 9'b110_000_101; // Magenta3
		8'ha4: color = 9'b110_000_110; // Magenta3
		8'ha5: color = 9'b110_000_111; // Magenta2
		8'ha6: color = 9'b110_010_000; // DarkOrange3
		8'ha7: color = 9'b110_010_010; // IndianRed
		8'ha8: color = 9'b110_010_100; // HotPink3
		8'ha9: color = 9'b110_010_101; // HotPink2
		8'haa: color = 9'b110_010_110; // Orchid
		8'hab: color = 9'b110_010_111; // MediumOrchid1
		8'hac: color = 9'b110_100_000; // Orange3
		8'had: color = 9'b110_100_010; // LightSalmon3
		8'hae: color = 9'b110_100_100; // LightPink3
		8'haf: color = 9'b110_100_101; // Pink3
		8'hb0: color = 9'b110_100_110; // Plum3
		8'hb1: color = 9'b110_100_111; // Violet
		8'hb2: color = 9'b110_101_000; // Gold3
		8'hb3: color = 9'b110_101_010; // LightGoldenrod3
		8'hb4: color = 9'b110_101_100; // Tan
		8'hb5: color = 9'b110_101_101; // MistyRose3
		8'hb6: color = 9'b110_101_110; // Thistle3
		8'hb7: color = 9'b110_101_111; // Plum2
		8'hb8: color = 9'b110_110_000; // Yellow3
		8'hb9: color = 9'b110_110_010; // Khaki3
		8'hba: color = 9'b110_110_100; // LightGoldenrod2
		8'hbb: color = 9'b110_110_101; // LightYellow3
		8'hbc: color = 9'b110_110_110; // Grey84
		8'hbd: color = 9'b110_110_111; // LightSteelBlue1
		8'hbe: color = 9'b110_111_000; // Yellow2
		8'hbf: color = 9'b110_111_010; // DarkOliveGreen1
		8'hc0: color = 9'b110_111_100; // DarkOliveGreen1
		8'hc1: color = 9'b110_111_101; // DarkSeaGreen1
		8'hc2: color = 9'b110_111_110; // Honeydew2
		8'hc3: color = 9'b110_111_111; // LightCyan1
		8'hc4: color = 9'b111_000_000; // Red1
		8'hc5: color = 9'b111_000_010; // DeepPink2
		8'hc6: color = 9'b111_000_100; // DeepPink1
		8'hc7: color = 9'b111_000_101; // DeepPink1
		8'hc8: color = 9'b111_000_110; // Magenta2
		8'hc9: color = 9'b111_000_111; // Magenta1
		8'hca: color = 9'b111_010_000; // OrangeRed1
		8'hcb: color = 9'b111_010_010; // IndianRed1
		8'hcc: color = 9'b111_010_100; // IndianRed1
		8'hcd: color = 9'b111_010_101; // HotPink
		8'hce: color = 9'b111_010_110; // HotPink
		8'hcf: color = 9'b111_010_111; // MediumOrchid1
		8'hd0: color = 9'b111_100_000; // DarkOrange
		8'hd1: color = 9'b111_100_010; // Salmon1
		8'hd2: color = 9'b111_100_100; // LightCoral
		8'hd3: color = 9'b111_100_101; // PaleVioletRed1
		8'hd4: color = 9'b111_100_110; // Orchid2
		8'hd5: color = 9'b111_100_111; // Orchid1
		8'hd6: color = 9'b111_101_000; // Orange1
		8'hd7: color = 9'b111_101_010; // SandyBrown
		8'hd8: color = 9'b111_101_100; // LightSalmon1
		8'hd9: color = 9'b111_101_101; // LightPink1
		8'hda: color = 9'b111_101_110; // Pink1
		8'hdb: color = 9'b111_101_111; // Plum1
		8'hdc: color = 9'b111_110_000; // Gold1
		8'hdd: color = 9'b111_110_010; // LightGoldenrod2
		8'hde: color = 9'b111_110_100; // LightGoldenrod2
		8'hdf: color = 9'b111_110_101; // NavajoWhite1
		8'he0: color = 9'b111_110_110; // MistyRose1
		8'he1: color = 9'b111_110_111; // Thistle1
		8'he2: color = 9'b111_111_000; // Yellow1
		8'he3: color = 9'b111_111_010; // LightGoldenrod1
		8'he4: color = 9'b111_111_100; // Khaki1
		8'he5: color = 9'b111_111_101; // Wheat1
		8'he6: color = 9'b111_111_110; // Cornsilk1
		8'he7: color = 9'b111_111_111; // Grey100
		8'he8: color = 9'b000_000_000; // Grey3
		8'he9: color = 9'b000_000_000; // Grey7
		8'hea: color = 9'b000_000_000; // Grey11
		8'heb: color = 9'b001_001_001; // Grey15
		8'hec: color = 9'b001_001_001; // Grey19
		8'hed: color = 9'b001_001_001; // Grey23
		8'hee: color = 9'b010_010_010; // Grey27
		8'hef: color = 9'b010_010_010; // Grey30
		8'hf0: color = 9'b010_010_010; // Grey35
		8'hf1: color = 9'b011_011_011; // Grey39
		8'hf2: color = 9'b011_011_011; // Grey42
		8'hf3: color = 9'b011_011_011; // Grey46
		8'hf4: color = 9'b100_100_100; // Grey50
		8'hf5: color = 9'b100_100_100; // Grey54
		8'hf6: color = 9'b100_100_100; // Grey58
		8'hf7: color = 9'b100_100_100; // Grey62
		8'hf8: color = 9'b101_101_101; // Grey66
		8'hf9: color = 9'b101_101_101; // Grey70
		8'hfa: color = 9'b101_101_101; // Grey74
		8'hfb: color = 9'b110_110_110; // Grey78
		8'hfc: color = 9'b110_110_110; // Grey82
		8'hfd: color = 9'b110_110_110; // Grey85
		8'hfe: color = 9'b111_111_111; // Grey89
		8'hff: color = 9'b111_111_111; // Grey93
		default: color = 9'b111_111_111;
	endcase
end

endmodule

module FontShapeRenderer (
    input clk,
    input rst,
    input [7:0] char,
    input []

);

parameter COLOR_NUMBERS = 4;

endmodule // FontShapeRender